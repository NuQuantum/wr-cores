library ieee;
use ieee.std_logic_1164.all;

package wr_txtsu_pkg is

-- t_txtsu_timestamp was here, but now it's moved to wr_endpoint_pkg.
  
end wr_txtsu_pkg;
